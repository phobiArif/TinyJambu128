library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

--PROGRAM de

entity de is
	port(
		clock : in std_logic;
		ne, ade, pe, sur, fb_en, pbade, pbce, sre, shift, cge, cgr, cre, re, te, tag1, tag2, mr, ps, mge : out std_logic;
		nscd, adscd, pscd, fbd, pbd, cgd, rd, td, pd : in std_logic;
		lim : out std_logic_vector(9 downto 0);
		cycle : in std_logic_vector(2 downto 0);
		fb : out std_logic_vector(2 downto 0);
		rx : in std_logic;
		mlen : in std_logic_vector(6 downto 0)
	);
end de;

architecture main of de is
	type keadaan is (
		idle, rxs, ks, fns, pn, usn,
		fads, pad, usad, pbad, fps,
		pp, usp, gm, pbp, fst1, fst2, pt1,
		pt2, gt1, gt2, tx
	);
	signal state : keadaan := idle;
begin
	process(all)
	begin
		if clock'event and clock = '1' then
			case state is
				when idle =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '1';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '0';
					shift <= '0';
					cge <= '0';
					cgr <= '1';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '1';
					ps <= '0';
					mge <= '0';
					if rx = '0' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '0';
						shift <= '0';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '1';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						ps <= '0';
						mge <= '0';
						state <= rxs;
					end if;
				when rxs =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '0';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '1';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					mge <= '0';
					if rd = '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '1';
						shift <= '1';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						ps <= '1';
						mge <= '0';
						lim <= conv_std_logic_vector(1023,10);
						state <= ks;
					end if;



					when fps =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '1';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					fb <= "101";
					mge <= '0';
					if fbd = '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '1';
						shift <= '1';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						ps <= '1';
						lim <= conv_std_logic_vector(1023,10);
						state <= pp;
						mge <= '0';
					end if;


					when pp =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '1';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '1';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '1';
					lim <= conv_std_logic_vector(1023,10);
					if pd <= '1' then
						ne <= '0';
						ade <= '0';
						pe <= '1';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '1';
						shift <= '0';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						ps <= '0';
						state <= usp;
						mge <= '0';
					end if;
				when usp =>
					ne <= '0';
					ade <= '0';
					pe <= '1';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '1';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					mge <= '1';
					if pscd = '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '1';
						shift <= '0';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						mge <= '0';
						ps <= '0';
						state <= usp;
					end if;
				when gm =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '1';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					mge <= '1';
					if cgd = '1' then
						if cycle < (mlen(6 downto 5)) + 1 then
							ne <= '0';
							ade <= '0';
							pe <= '0';
							sur <= '0';
							fb_en <= '1';
							pbade <= '0';
							pbce <= '0';
							sre <= '1';
							shift <= '0';
							cge <= '0';
							cgr <= '0';
							cre <= '0';
							re <= '0';
							te <= '0';
							tag1 <= '0';
							tag2 <= '0';
							mr <= '0';
							ps <= '0';
							state <= fps;
							fb <= "101";
							mge <= '0';
						else
							if mlen(4 downto 0) = 0 then
								ne <= '0';
								ade <= '0';
								pe <= '0';
								sur <= '1';
								fb_en <= '1';
								pbade <= '0';
								pbce <= '0';
								sre <= '1';
								shift <= '0';
								cge <= '0';
								cgr <= '0';
								cre <= '0';
								re <= '0';
								te <= '0';
								tag1 <= '0';
								tag2 <= '0';
								mr <= '0';
								ps <= '0';
								state <= fst1;
								fb <= "111";
								mge <= '1';
							else
								ne <= '0';
								ade <= '0';
								pe <= '0';
								sur <= '0';
								fb_en <= '0';
								pbade <= '0';
								pbce <= '1';
								sre <= '1';
								shift <= '0';
								cge <= '0';
								cgr <= '0';
								cre <= '0';
								re <= '0';
								te <= '0';
								tag1 <= '0';
								tag2 <= '0';
								mr <= '0';
								ps <= '0';
								state <= pbp;
								mge <= '0';
							end if;
						end if;
					end if;
				when pbp =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '1';
					sre <= '1';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					mge <= '1';
					if pbd = '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '1';
						pbade <= '0';
						pbce <= '0';
						sre <= '1';
						shift <= '0';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						ps <= '0';
						state <= fst1;
						fb <= "111";
						mge <= '1';
					end if;
				when fst1 =>				
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '1';
					fb_en <= '1';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					fb <= "111";
					mge <= '1';
					if fbd = '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '1';
						shift <= '1';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						ps <= '1';
						lim <= conv_std_logic_vector(1023,10);
						state <= pt1;
						mge <= '1';
					end if;
				when pt1 =>	
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '1';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '1';
					lim <= conv_std_logic_vector(1023,10);
					mge <= '1';
					if pd = '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '0';
						shift <= '0';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '1';
						tag2 <= '0';
						mr <= '0';
						ps <= '0';
						state <= gt1;
						mge <= '1';
					end if;
				when gt1 =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '1';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					state <= fst2;
					fb <= "111";
					mge <= '1';
				when fst2 =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '1';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					fb <= "111";
					mge <= '1';
					if fbd <= '1' then	
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '1';
						shift <= '1';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '0';
						ps <= '1';
						lim <= conv_std_logic_vector(639,10);
						state <= pt2;
						mge <= '1';
					end if;
				when pt2 =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '1';
					shift <= '1';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '0';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '1';
					lim <= conv_std_logic_vector(639,10);
					mge <= '1';
					if pd <= '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '0';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '0';
						shift <= '0';
						cge <= '0';
						cgr <= '0';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '1';
						mr <= '0';
						ps <= '0';
						state <= gt2;
						mge <= '1';
					end if;
				when gt2 =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '0';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '1';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					state <= tx;
					mge <= '1';
				when tx =>
					ne <= '0';
					ade <= '0';
					pe <= '0';
					sur <= '0';
					fb_en <= '0';
					pbade <= '0';
					pbce <= '0';
					sre <= '0';
					shift <= '0';
					cge <= '0';
					cgr <= '0';
					cre <= '0';
					re <= '0';
					te <= '1';
					tag1 <= '0';
					tag2 <= '0';
					mr <= '0';
					ps <= '0';
					mge <= '1';
					if td = '1' then
						ne <= '0';
						ade <= '0';
						pe <= '0';
						sur <= '1';
						fb_en <= '0';
						pbade <= '0';
						pbce <= '0';
						sre <= '0';
						shift <= '0';
						cge <= '0';
						cgr <= '1';
						cre <= '0';
						re <= '0';
						te <= '0';
						tag1 <= '0';
						tag2 <= '0';
						mr <= '1';
						ps <= '0';
						state <= idle;
						mge <= '1';
					end if;
			end case;
		end if;
	end process;
end main;